`ifndef COMMON_VH
`define COMMON_VH

`define DIR_DOWN    0
`define DIR_UP      1

`define SHIFT_DIR_LEFT    0
`define SHIFT_DIR_RIGHT   1

`endif
