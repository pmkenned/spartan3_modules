`default_nettype none
`timescale 1ns / 1ps

module top(
    input wire clk,
    input wire [7:0] switches,
    input wire [3:0] buttons,
    output wire [7:0] leds,
    output wire [6:0] ss_abcdefg_l,
    output wire ss_dp_l,
    output wire [3:0] ss_sel_l
);

    wire rst;
    assign rst = buttons[3];

    assign leds[7:0] = 'b0;

    wire [31:0] bram_data_out;
    wire [3:0] bram_parity_out;
    wire [31:0] bram_data_in;
    wire [3:0] bram_parity_in;
    wire [8:0] bram_addr;
    wire bram_en;
    wire bram_ssr;
    wire bram_we;

    assign bram_data_in = 'b0;
    assign bram_parity_in = 'b0;
    assign bram_addr = {1'b0, switches};
    assign bram_en = 1'b1;
    assign bram_ssr = 1'b0;
    assign bram_we = 1'b0;

    ss_driver primary_ss_driver(
        .clk(clk),
        .rst(rst),
        .hex_digits(bram_data_out[15:0]),
        .ss_abcdefg_l(ss_abcdefg_l),
        .ss_dp_l(ss_dp_l),
        .ss_sel_l(ss_sel_l)
    );

    // RAMB16_S36: 512 x 32 + 4 Parity bits Single-Port RAM
    RAMB16_S36 #(
        .INIT(36'h000000000),  // Value of output RAM registers at startup
        .SRVAL(36'h000000000), // Output value upon SSR assertion
        .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

        // The following INIT_xx declarations specify the initial contents of the RAM
        // Address 0 to 127
        .INIT_00(256'h00112233_44556677_8899aabb_ccddeeff_feedbabe_deadbeef_01234567_89abcdef),
        .INIT_01(256'haaaaaaaa_bbbbbbbb_cccccccc_dddddddd_eeeeeeee_ffffffff_11111111_22222222),
        .INIT_02(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_03(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_04(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_05(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_06(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_07(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_08(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_09(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_0A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_0B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_0C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_0D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_0E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_0F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        // Address 128 to 255
        .INIT_10(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_11(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_12(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_13(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_14(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_15(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_16(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_17(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_18(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_19(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_1A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_1B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_1C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_1D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_1E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_1F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        // Address 256 to 383
        .INIT_20(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_21(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_22(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_23(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_24(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_25(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_26(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_27(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_28(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_29(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_2A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_2B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_2C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_2D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_2E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_2F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        // Address 384 to 511
        .INIT_30(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_31(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_32(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_33(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_34(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_35(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_36(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_37(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_38(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_39(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_3A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_3B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_3C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_3D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_3E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
        .INIT_3F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),

        // The next set of INITP_xx are for the parity bits
        // Address 0 to 127
        .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
        // Address 128 to 255
        .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
        // Address 256 to 383
        .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
        // Address 384 to 511
        .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
        .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
    ) RAMB16_S36_inst (
        .DO(bram_data_out),
        .DOP(bram_parity_out),
        .ADDR(bram_addr),
        .CLK(clk),
        .DI(bram_data_in),
        .DIP(bram_parity_in),
        .EN(bram_en),
        .SSR(bram_ssr),
        .WE(bram_we)
    );

endmodule

module hex_to_ss
#(parameter ROTATE=0)
(
    input wire [3:0] hex,
    output reg [6:0] ss_abcdefg_l
);

    always @(hex) begin
        case (hex)
            4'h0: ss_abcdefg_l = ROTATE ? 7'b0000001 : 7'b0000001;
            4'h1: ss_abcdefg_l = ROTATE ? 7'b1111001 : 7'b1001111;
            4'h2: ss_abcdefg_l = ROTATE ? 7'b0010010 : 7'b0010010;
            4'h3: ss_abcdefg_l = ROTATE ? 7'b0110000 : 7'b0000110;
            4'h4: ss_abcdefg_l = ROTATE ? 7'b1101000 : 7'b1001100;
            4'h5: ss_abcdefg_l = ROTATE ? 7'b0100100 : 7'b0100100;
            4'h6: ss_abcdefg_l = ROTATE ? 7'b0000100 : 7'b0100000;
            4'h7: ss_abcdefg_l = ROTATE ? 7'b1110001 : 7'b0001111;
            4'h8: ss_abcdefg_l = ROTATE ? 7'b0000000 : 7'b0000000;
            4'h9: ss_abcdefg_l = ROTATE ? 7'b1100000 : 7'b0001100;
            4'ha: ss_abcdefg_l = ROTATE ? 7'b1000000 : 7'b0001000;
            4'hb: ss_abcdefg_l = ROTATE ? 7'b0001100 : 7'b1100000;
            4'hc: ss_abcdefg_l = ROTATE ? 7'b0000111 : 7'b0110001;
            4'hd: ss_abcdefg_l = ROTATE ? 7'b0011000 : 7'b1000010;
            4'he: ss_abcdefg_l = ROTATE ? 7'b0000110 : 7'b0110000;
            4'hf: ss_abcdefg_l = ROTATE ? 7'b1000110 : 7'b0111000;
            default: ss_abcdefg_l = 7'b1111111;
        endcase
    end

endmodule

module ss_driver
#(parameter ROTATE = 0)
(
    input wire clk,
    input wire rst,
    input wire [15:0] hex_digits,
    output reg [6:0] ss_abcdefg_l,
    output wire ss_dp_l,
    output wire [3:0] ss_sel_l
);

    reg [19:0] clk_cnt;
    wire clk_191Hz;
    assign clk_191Hz = clk_cnt[17];

    always @(posedge clk, posedge rst) begin
        if (rst) begin
            clk_cnt <= 20'b0;
        end else begin
            clk_cnt <= clk_cnt + 20'b1;
        end
    end

    reg [3:0] cycler;
    wire [3:0] cycler_n;
    wire [6:0] ss_array_l [3:0];

    assign cycler_n[1] = cycler[0];
    assign cycler_n[2] = cycler[1];
    assign cycler_n[3] = cycler[2];
    assign cycler_n[0] = cycler[3];

    assign ss_sel_l = ~cycler;

    always @(posedge clk_191Hz, posedge rst) begin
        if (rst) begin
            cycler <= 4'b1;
        end else begin
            cycler <= cycler_n;
        end
    end

    always @(cycler, ss_array_l[0], ss_array_l[1], ss_array_l[2], ss_array_l[3]) begin
        case (cycler)
            4'b0001: ss_abcdefg_l = ss_array_l[0];
            4'b0010: ss_abcdefg_l = ss_array_l[1];
            4'b0100: ss_abcdefg_l = ss_array_l[2];
            4'b1000: ss_abcdefg_l = ss_array_l[3];
            default: ss_abcdefg_l = 7'b1111111;
        endcase
    end

    assign ss_dp_l = 1'b1;

    hex_to_ss #(.ROTATE(ROTATE)) hts0(.hex(hex_digits[3:0]),   .ss_abcdefg_l(ss_array_l[0]));
    hex_to_ss #(.ROTATE(ROTATE)) hts1(.hex(hex_digits[7:4]),   .ss_abcdefg_l(ss_array_l[1]));
    hex_to_ss #(.ROTATE(ROTATE)) hts2(.hex(hex_digits[11:8]),  .ss_abcdefg_l(ss_array_l[2]));
    hex_to_ss #(.ROTATE(ROTATE)) hts3(.hex(hex_digits[15:12]), .ss_abcdefg_l(ss_array_l[3]));

endmodule
